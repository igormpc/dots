BZh91AY&SYH�Y N_�Py���߰����P��$*�H���	���dɓ#	�i�F& ��A�ɓ&F�L�LD@SDS�l��jc&�A��d�4f�9�14L�2da0M4����$AM4i0��S�S�=Q�4 �<���M�
�$,&$���"�ȣ����b�blؓG�+4�v21(1��E�;�����Ζ�UGS������
?�tP�LJ+�����fT�p$���3Ы���᱐sp�B�Hrnj3����j�Zv��'�d�,�`�1yuXU��� �ؐ�6�UuFs�4yns�5�J�F��mgmF�R���^/ŽxʷP�Z2�)���.ՔND��I��4s�ʰ�aå2E�{M�W1bL1��/��C��#����A�*�h��/n�myXH��SM�G�qc���m���� t#����J�^%�+�1\���;�.�K
+�b��&����I�(�P�2C���u��Q)�Ƙ<�e�Z�1a`�F�֛�­,�Sg'�f��K�v{t^���=��l���}�)c6�spF��E�P�ߊ^���3�XC���N`�],���r���zK<s�7��i�}�gD���D��?�5#�p�ψ��Q)6>f����Z~���R�S�������o��8)J�\��=amt'�/��Q{K�G����-]X���ө0�@sծ�R*ƃ�Zx����d���.q�X!��T��hA`p^^a���͂LZ!�xE�ER����{��NqsHzѦ��9�d�th���Α������.�P��J��Z�h�G�e�F�n�9��<*`k�����{�ˀ��g<��o�d���:S�:��[T娻�7
�t�|�ǙRp��X[&7��jz���)�v��p)R72��/&��i�C���Q�x%�*V�VJX�5�w`J0�g�L�Ԝ׃Y3�ΊJM/u@:�\!��̕`!N�r^�Rڙ���9��ȏ�_�Z�*l&<�nv��=OC�M�����9$pN��\�:NNS��$��GDR�u���V�Ve)ӥo땰��~I�8͟�B4GnFP�X�������G������Y�')Q&-��[cdi����V��jvm8�S{&�tbJ;0�Ӊ�����X]8��${����Cq�l�s�LLh�G,c�G�NiU)S���J�Ѵ3?���)�G}j�